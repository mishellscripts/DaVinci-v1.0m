// Name: alu.v
// Module: ALU
// Input: OP1[32] - operand 1
//        OP2[32] - operand 2
//        OPRN[6] - operation code
// Output: OUT[32] - output result for the operation
//
// Notes: 32 bit combinatorial ALU
// 
// Supports the following functions
//	- Integer add (0x1), sub(0x2), mul(0x3)
//	- Integer shift_rigth (0x4), shift_left (0x5)
//	- Bitwise and (0x6), or (0x7), nor (0x8)
//  - set less than (0x9)
//
// Revision History:
//
// Version	Date		Who		email			note
//------------------------------------------------------------------------------------------
//  1.0     Sep 10, 2014	Kaushik Patra	kpatra@sjsu.edu		Initial creation
//  1.1     Oct 19, 2014        Kaushik Patra   kpatra@sjsu.edu         Added ZERO status output
//------------------------------------------------------------------------------------------
//
`include "prj_definition.v"
module ALU(OUT, ZERO, OP1, OP2, OPRN);
// input list
input [`DATA_INDEX_LIMIT:0] OP1; // operand 1
input [`DATA_INDEX_LIMIT:0] OP2; // operand 2
input [`ALU_OPRN_INDEX_LIMIT:0] OPRN; // operation code

// output list
output [`DATA_INDEX_LIMIT:0] OUT; // result of the operation.
output ZERO; // zero flag

// simulator internal storage - this is not h/w register
reg [`DATA_INDEX_LIMIT:0] result;
reg [`DATA_INDEX_LIMIT:0] zero;

// whenever op1, op2, or oprn changes
always @(OP1 or OP2 or OPRN)
begin
    case (OPRN)
	`ALU_OPRN_WIDTH'h01 : result = OP1 + OP2; // addition
	`ALU_OPRN_WIDTH'h02 : result = OP1 - OP2; // subtraction
	`ALU_OPRN_WIDTH'h03 : result = OP1 * OP2; // multiplication
	`ALU_OPRN_WIDTH'h04 : result = OP1 >> OP2; // shift right
	`ALU_OPRN_WIDTH'h05 : result = OP1 << OP2; // shift left
	`ALU_OPRN_WIDTH'h06 : result = OP1 & OP2; // bitwise and
	`ALU_OPRN_WIDTH'h07 : result = OP1 | OP2; // bitwise or
	`ALU_OPRN_WIDTH'h08 : result = ~(OP1 | OP2); // bitwise nor
	`ALU_OPRN_WIDTH'h09 : result = (OP1 < OP2)?1:0;// set less than
        default: result = `DATA_WIDTH'hxxxxxxxx;            
    endcase
    if (result === 0)
       zero = 1'b1;
    else
       zero = 1'b0;
end

assign OUT = result;
assign ZERO = zero;

endmodule
